----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:39:25 07/31/2009 
-- Design Name: 
-- Module Name:    top - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity top is
	port ( sys_clk: in std_logic;
			 Led: out std_logic_vector(7 downto 0));
end top;

architecture Behavioral of top is
	signal CAPTURE: std_logic;
	signal UPDATE: std_logic;
	signal UPDATE_sync: std_logic;
	signal DRCK1: std_logic;
	signal last_DRCK1: std_logic;
	signal TDI: std_logic;
	signal TDO1: std_logic;
	signal SEL1: std_logic;
	signal SEL1_sync: std_logic;
	signal SHIFT: std_logic;
	signal RESET: std_logic;
	signal ctl: std_logic_vector(7 downto 0);
	signal addr: std_logic_vector(15 downto 0);
	signal data_wr: std_logic_vector(15 downto 0);
	signal data_rd: std_logic_vector(15 downto 0);
	signal shift_in: std_logic_vector(39 downto 0);
	signal shift_out: std_logic_vector(39 downto 0);
	signal ram_we: std_logic := '0';
	signal last_update: std_logic;
begin
	JTAG : BSCAN_SPARTAN3
       port map (CAPTURE => CAPTURE,
                 DRCK1 => DRCK1,
                 DRCK2 => open,
                 RESET => RESET,
                 SEL1 => SEL1,
                 SEL2 => open,
                 SHIFT => SHIFT,
                 TDI => TDI,
                 UPDATE => UPDATE,
                 TDO1 => TDO1,
                 TDO2 => open); 

   RAMB16_S18_S18_inst : RAMB16_S18_S18
   generic map (
      INIT_A => X"00000", --  Value of output RAM registers on Port A at startup
      INIT_B => X"00000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"00000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"00000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
      -- The follosing INIT_xx declarations specify the intiial contents of the RAM
      -- Address 0 to 255
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 256 to 511
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 512 to 767
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 768 to 1023
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Address 0 to 255
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 256 to 511
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 512 to 767
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 768 to 1023
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => data_rd,      -- Port A 16-bit Data Output
      DOB => open,      -- Port B 16-bit Data Output
      DOPA => open,    -- Port A 2-bit Parity Output
      DOPB => open,    -- Port B 2-bit Parity Output
      ADDRA => addr(9 downto 0),  -- Port A 10-bit Address Input
      ADDRB => "0000000000",  -- Port B 10-bit Address Input
      CLKA => sys_clk,    -- Port A Clock
      CLKB => sys_clk,    -- Port B Clock
      DIA => data_wr,      -- Port A 16-bit Data Input
      DIB => x"0000",      -- Port B 16-bit Data Input
      DIPA => "00",    -- Port A 2-bit parity Input
      DIPB => "00",    -- Port-B 2-bit parity Input
      ENA => '1',      -- Port A RAM Enable Input
      ENB => '0',      -- PortB RAM Enable Input
      SSRA => '0',    -- Port A Synchronous Set/Reset Input
      SSRB => '0',    -- Port B Synchronous Set/Reset Input
      WEA => ram_we,      -- Port A Write Enable Input
      WEB => '0'       -- Port B Write Enable Input
   );

	process(sys_clk)
	begin
	
		if rising_edge(sys_clk) then
		
			ram_we <= '0';
			
			--last_DRCK1 <= DRCK1;
			SEL1_sync <= SEL1;
			
			UPDATE_sync <= UPDATE;
			last_update <= UPDATE_sync;
			
			if last_update = '0' and UPDATE_sync = '1' and SEL1_sync = '1' then
				ctl <= shift_in(39 downto 32);
				addr <= shift_in(31 downto 16);
				data_wr <= shift_in(15 downto 0);
				ram_we <= shift_in(32);
				Led <= shift_in(39 downto 32);			
			end if;
			
		end if;
	end process;
			
	process(DRCK1)
	begin
	
		if rising_edge(DRCK1) then
			
			if SEL1 = '1' then
			
				if SHIFT = '1' then
					shift_in <= shift_in(38 downto 0) & TDI;
					shift_out <= shift_out(38 downto 0) & '0';
				else
					shift_out <= ctl & addr & data_rd;
				end if;
			
			end if;
			
			--if SEL1 = '1' and SHIFT = '1' then
				--shift_in <= shift_in(38 downto 0) & TDI;
				--shift_out <= shift_out(38 downto 0) & '0';
			--end if;
			
			--if SEL1 = '1' and CAPTURE = '1' then
				--shift_out <= ctl & addr & data_rd;
			--end if;
			
		end if;
	
	end process;

	--process(DRCK1)
	--begin
	
--		if falling_edge(DRCK1) and SHIFT='1' and SEL1='1' then
	--		shift_out <= shift_out(38 downto 0) & '0';
		--	TDO1 <= shift_out(38);
		--end if;
	
	--end process;

	TDO1 <= shift_out(39);

end Behavioral;

